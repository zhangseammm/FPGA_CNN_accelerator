module tb_module_quan(

   );
endmodule